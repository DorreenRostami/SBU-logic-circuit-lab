`timescale 1ns / 1ps
module xor_gate(
    input A,
    input B,
    output C
    );

	assign C = A ^ B;
endmodule
