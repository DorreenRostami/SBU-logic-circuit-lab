`timescale 1ns / 1ps
module not_gate(
    input A,
    output B
    );

	assign B = ~A;
endmodule
